`ifndef __param_ram__
`define __param_ram__

`define DWIDTH 32
`define AWIDTH 32
`define LWIDTH 2
`define  WORDS 16384

`endif