`ifndef __param_csr_addr__
`define __param_csr_addr__


`define CSR_ADDR_MTVEC 12'h305
`define CSR_ADDR_MEPC 12'h341
`define CSR_ADDR_MCAUSE 12'h342
`define CSR_ADDR_NONE 12'hfff

`endif
