`ifndef __param_pc_mux__
`define __param_pc_mux__

`define SEL_PC_WIDTH 2

`define SEL_PC_NONE 2'b00
`define SEL_PC_ADD4 2'b01
`define SEL_PC_JAL 2'b10
`define SEL_PC_JALR 2'b11

`endif
