`ifndef __param_pc_mux__
`define __param_pc_mux__

`define PC_SEL_WIDTH 2
`define PC_SEL_NONE 2'b00
`define PC_SEL_ADD4 2'b01
`define PC_SEL_JAL 2'b10
`define PC_SEL_JALR 2'b11

`endif
