`ifndef __param_src_a_mux__
`define __param_src_a_mux__


`define SEL_SRC_A_WIDTH 2

`define SEL_SRC_A_PC  2'h1
`define SEL_SRC_A_RS1 2'h2
`define SEL_SRC_A_IMM 2'h3


`endif
